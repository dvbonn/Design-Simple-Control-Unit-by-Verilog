library verilog;
use verilog.vl_types.all;
entity MIPSCPU_tb is
end MIPSCPU_tb;
